bind fifo fifo_checker_sva check_fifo(clk, rst, rqst_i, gnt_o);
